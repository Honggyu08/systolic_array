module PE(clk, inp, add, outp);

input clk;
input inp;
input add;

output outp;


